
interface intf();
    // ------------------- port declaration-------------------------------------
    logic [7:0] in;
    logic [8:0] out;
    //--------------------------------------------------------------------------    
endinterface


module bin2ex3(in,out);
    input  [7:0]  in;
    output [8:0] out;

    assign out=in+3;

endmodule